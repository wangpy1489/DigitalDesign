library verilog;
use verilog.vl_types.all;
entity pipe_computer_sim is
end pipe_computer_sim;
